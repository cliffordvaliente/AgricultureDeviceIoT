PK   �WW��?�(  �    cirkitFile.json�k��F������Z,d$�����e��cÞ�@��[�r�_�z<����fPU]*&)%'l�^�K$���<$3��j_���_ov�n��n���ݯ^Qv�zW�۟��O�����~}ح���߭^��'���f��m��۬]Uo:��*�,q}�&�5�[�iY���~m�f����7�+�X��I� U0k+f�*�u*f�*��3H�:3H�:3H̺3H̺3H̺3H|��J��� �Jy�$y�Kx
y�Kx
y�Kx
y�Kx
y�Kx
y�Kx
y�Kx
y�K����v�%<��v�%<`�)��V^;��B^;��B^;��B^;��B^;��B^;��B^;���k�X�S�k�X�S�k�X�S l��v���)����)����)����)����)����)�0k'��b	O!��b	O!��b	O!��b	O��)��N^;��B^;��B^;��B^;��B^;�f��k�X�S�k�X�S�k�X�S�k�X�S�k�X�S n�kg&��b	O!��b	O!��b	O!��b	���S,�)�S,�)�3�x����'�z{�������o��? ���r�=�mv?���w��u�5٦�7I��*qY[%%�}�7iQe6�2S��
Fr�aW�d"�Y�{��{JGX:����Yl���kL�lSPRP_$κ4���I\�6�����fM�l��0�N�aO�a��QHw�^��J�awذtSq�ޫ�&i]���.)�.O�uM^���fm���a~��{�;��B�����f��6�96��d�L�W�+[�^��&iL]$�9�Q]U.�v�3��v(a�̺�Ʈ��JG!��G@*�6�6�P:���Ӟ`�v�X>��s���������-�=���|�l08~`3��#0?���Ua����c���GX>������}���|�<8~`Â�#0?��ش`�������,��x��>�`���s=���,��x�
8~�{H`�����5�������|<3?�������4���X>��l,p����G`>�G��`���3����,��x�8~`���	���NmQ�uS�IZ6i�6E�Ԏ��,˞�Ҧ��1��<a�غ�|W�J�����,Mp����G|W�Jك�<5z�a����'Ղ�~z���0�`Ô����|<�?�a�����`��6LX>���qp���	�G`>����0a������&,���� 6~�z�|��&	�������|��?������S���X>�qKp���p�����@���,����	8~`���#07`��?�|���1�������|��?��������`㗁����|�h?������[$���X>�qs'p����G`>nK��`������C��GO����?2�����������X>�q�5p����G`>n��`���-������G`>n����|�?5'mR��mܢ{�w�������e���=~N����2.�	BT�C�$_=nn��K�,����4IT7#�a%�f����Qd/;I�7�:��p�q�ץ��l�q���]Pe{���CdT�0�}�n>n�p�r�6D�̳��]�|sdI�B�CPx��\���(^k�t�q����S>x	�����̗n?��Q#�T��v�\��sc¸���y�Y��p�`P��D��${MTe�W^�"Duvx����-�܉-�e1�����K��?�#{!��U.�9���d1#��a����o�/��3N�����a�N�����XrIb�9v|5�Y��y��@�\�;�Ǝ�_=?r��|~�����5j���s�$q�E���:`!�n�?W�c���$=�Ƿ&$,��5�K�o`և�z����W�~~�_�2%h��d����%d���!	>ob�@B�O�"���,�$d�d�!	>c�@B�O�"����$dx��!	�a<*����+۰�M�R2ø���+�(%3��@L��M��R2�-�������p����V�QJf�Yb�qpX��:�R2Í"��[XG)����	V�-�����p+
���V�QJf�u��:���8J�;pWRp�R`u<��q�w��1��x
��(%�c���V�QJ�����V�QJ�u
���V�QJ�	Ƅ�&��(��V�QJ����V�QJ�����V�QJ�iv�V�3XG)qG��g�:�R��0&��M��MX�`u�ĳ�aL�:���8J�g�Ø`u<��q�ς�1��x��sJ�g,�'��U�i��`r�W��K��#+�էv��'�c�:�����+����]�*0�!+"_5X�z���
��k0T�Ϳ0q� �D dE��Y����U�q�`���u�,�q�0LBVD�j�����\WVRa5�qs1�*0��AP7��u�zVRa�g�u����R�%Z~�Y'�J�K�v��.�1^��ThI���5׉���R�%Z~f^'�:L��th�����0Zҡ�9:��qb*��C�s1tb���ThI�����VǑ�В-ύщ��+S�%Z��scAǗ�В-�U҉��/S�%Z�s�[�;b:�L�����VǗ�В-ρӉ��/S�%Z�˧[_�BK:�<'Q'�:�L��thyn�Nlu|�
-���Q����2Zҡ5/�P"c���Th�V����㶚��t|�-�Z�c&2�:�L�6l��[_���2Zҡ��:�UzZQ�qE_����TǗ�В-��׉��/S�%Z�1�[_�BK:��+A'�:�L��th��Nlu|�
-��r�
����2Zҡ�*�u:�L��th���Nlu|�
-��rO����2Zҡ��.:���e*��C�=jtb�4�LǗ��r�����2Zҡ�A:���e*��C˽�tb���ThI��{8��VǗ�В-��҉��/S�%Z�LǗ�В-�Ӊ��/S�%Z�q�[_�BK:�ܫM'�:�L��th��Nlu|�
-��r�<��*u�Pj���2_���2Zҡ�^�:���e*��C�=ub���ThI��{K��VǗ�В-��T�m���ThI���V�E�6������e��/�-[_6A>#����Δyչ"�e�Uk���E�����uQ���0�;~��coڬO+��L7م*饸4�u�)()�/g]�T}�$�jWQ�V}s�K�Sv��({�E�$}���B��.�K_�Q��ؾP�]�GQ*d��1_�2�y|���+���X�Ju�8��:P�b�w���Ke0�;�ݥ23}���`Rx��Kef�/��8�K�o$U�1�뮐soJ]*�����.�q��q2�Y\�M&�����l��cS�$g�X��T�7�Z��֒�.�Ͻ'�d���~<욤um�GD�Kʾ�k]��iG}���ƨ�űt���tƌR�x<�E��M�&i٤��]R;�1.˞�ҦUǸ��EQ*ǯQ*��1��^��Q*��R!�R�x��R�x��R�x��R�y��Ҭ3��o�]��q2�R���I/U�8��v%N�ԯ�2���á>t�W??�.�����a_ߝ.�H�UB2CE����P]!D !3TjH�UB2�B2��B2ÙB2�YB2�3.�D�6�l��6�
7J�&X�&X�F)�����+�(%s��a��p�q��9^�0�긅�q��9^��0��߸8��[XG)��UY��[XG)���b��[XG)��l��[XG)��5v����V�QJ܇Ƅ�������)�����_�	V�SXG)q"����:�R�~80&Xw�:�R��+0&Xw�:�R�~0&�5q�EqXw�:�R�0&Xw�:�R�> 0&Xw�:�R�y�[?�:���8J��9Ø`u<��q�ϫ�1��n�no��x��(%��c���V�QJ<����9����x~�	V�sX�SZ>W+��V=N���
+���u0�
��+���u0�
��+���uЗ�
��+��zߥנ%$�����A*qڱ@"��J*�~��נ$���j�A�*0����j�A�*0����j�A��*0�������ǥBK:��l�Nl�\�����]�c�H�y�В-?k�[��BK:��̼Nlu�
-����:��qa*��C�stb���ThI���b��VǍ�В-�)щ��#S�%Z��[W�BK:�<�G�Ƃ�/S�%Z���[_�BK:�<�J'�JwĔn���2��ˬ�/S�%Z��[_�BK:�<�O'�:�L��thyN�Nlu|�
-����J����2Zҡ�9�:���e*��C�s]ub���ThI�����<����ThI�����VǗ�В-ϡ։��/S�%Z��[���W��e��/Ku|�
-����|����2Zҡ�:���e*��C˽tb���ThI��{>��VǗ�В-��Љ��/S�%Z���[���ThI��{���VǗ�В-�Dщ��/S�%Z��[_�BK:�ܣF'�J3ɔ����2��˜�/S�%Z��[_�BK:���H'�:�L��th���Nlu|�
-��r/*����2Zҡ�Z*��t|�
-��ro0����2Zҡ�g:���e*��C˽�tb���ThI��{���VǗ�В-��Ӊ�R��6:�,��e��/S�%Z�e�[_�BK:�ܓQ'�:�L��th���Nlu|�
-��r�L���:�L��th�קNlu|�
-��r�R����2Z��=y!�)�sEb�ޫ6�$���dc3�?�����üPe�7�B��n�Uf�x?�4�u�)()�/g]�T}�$�jWQ�V}s9.Q*��r1.y�d�*�$yc��em����IߤE��<�L}�E�\�EQ*�_tqOG���X_�2�}��L�*3�����
_�2��{iց���s��]*��߹��.��d�ܫj��`rxKe0Y<��ե2������.��d��[?��`�x�ݚKe0Y<�˥g]LϽ'�d���~<욤um�GD�Kʾ�k]��iG}���ƨ`X.�_cT.OmQ�uS�IZ6i�6E�Ԏ|�˲���iF��D�\�K��ŸD�`�r��D�\�2Q*�L����r��D�\�0qYJ^L�^���`���h/N�4�������z�������_�WdoV?m�����]�����~�۷�~����VKt�ct5����$��/�̐D^h�X4I*���o&Y�mTD^Z��Qy9��=�������.&V2�u��W����RU~t��`������+")�r0�L	�h/b�@��|D,�$O+�w�
���;�]}�d�`s�w�B���ZX��-�D{@8^��F�a�M�W�и׍%���ž}�9����?�ѩ��)������#���@�� �G)�B���Dh�� ���@`sv��hr �U�I��8�n��#�/ȿ�u<�k8H9�Hʁ�~�,�oc+Hhw	@��L ��k��� u�r���}(`���H�J�hs*'{Tv������߭��[���������n�aۮ^���e;��f�׍}"�o��Oy�J�\��)�fxnAH!�0�sB
����R�%��܅�B,a��6�b	3<�!�K��!�X�ϝ)���܊�l!�'�|�'
�\���r j(��\���r �(
�\�6�r j)��\�w�r ��S��9>p/�@�GR@=��z*�0�9R@=��z*�0�YR@=��z*�0�yR@=��z*�0ǙR+	��)���5�-6 ��GX|@=M�T��op �i
��r~C�POS@=�k� �z� �T����z� �T�����k�����z� �T��ݲ�z� �T��]��z� �T���}���4�S�w�p �i��r�F
�@܅B܆��PO��������5�� �POs@=�kp; ���zj,�:t5������Vf�&���j2렯�0�ACCat�|�3����z��|��>��5렍<NN,_0�"�=����x�8�A�x���F?_��7׬�f�8=H8�|���`�䲟��3h/�����W0yHv-�qz�pb��g�A�w�$~X�`��8�I4p5�ӻ0�A�w��������D���LHhB~�C�����!��!������E�ml���&���1D�0!�	�Yft�LHhB~C�o���!G�mV���&����1D0!�	��}t�.LHhB�w����)`BB�	t�>LHhB�!�^ڧ�	y�
:�h�&$4!ϳA��S���&�9B��}
��Є<�	C�O���f�c��)`BB�2t�>LHhB�&�h�&�?��JY�ݜ䏚�mKH8����3ؼh�	)�ŀ	��W�}d���hS��M��Є<aC�Se���Ц&E��mj���&䉺��M��Є<�C����'H�c�65`BB��ntѦLHhB����!�Ԁ		Mȓ��1th&$4!7@�m[���&�f��}
��Є܈C�O���H�c���)`Bn���!ڧ�		M��;�1D�0!�	��:�h�&$4!7MA��S���&�/��}
��Єܬ��S���&�F;��}
��Є�$C�O���c��)`BBrs&t�>LHhBn,��!|>>|B>ڧdh���}
��Є��C�O�����c��)`BBr#5t�>LHhBn�a��)`BB��ͦPAL�ѓu�wi��͋��bB��-`���>�y�k���7�Y�
�@��M���|/��/�����e��&�5����ޟo����Aϥoenf�Gm4^���)y�q�I^���]�}�6w�烟S��#+.���+�����K����o�@�jz��4I×�-�2/�t� ����)Ċ^P.���<_ȶT`��Όb����%�ix��H/�����M�a)&�y߆)O����o�Z*p&ǻ���g�$�ks?2]R�]�X뚼L;���԰m&�Qrö�|����ͤk�ܙ�1��a�h�h���E3�"J.�ܱ%����%V2;3Ƌ��ܹ"J���8j�3'��Ϝ����l�4'R{���ӛ�홺�7��3�<No����8�0�I��4q���/7�g�m�>���V�~^�X�ի�W|�q�p����*�>���osn
��fŻ�ӀS�kWO.yÕ��Z��aW�wH�!�Z6�ۡH�h� �qoy�[X���������-R�/=~��b2X1�����U6�t}�K��}��I٥mb�#OR�C�y/�?[[QR5��!E�&M�����.�;�s����զ��&�����")7U��uuc�ژ����Mi��$i�w���6i�"O�ޑ��g
~��i:�y[&��Y����wu�Ro���9}�~8��}w�]?n?��!��҄���yG8a���5��J�f��W�B�t&���(R��nt8����n�f�"G����.E.��	wkv)r�Nr����)�`���.�4��F�T������y'CW^H*�+��#9��o���\�7IC���@�8]t�&ę+��6Dt1*ę+��.Kt�-ę+�&Rt)1ę+��CDJC��zy�H6��.����y)J6��4l�s>�R��.EH#��9n҉
��r��?{�C�����n�;�jf�o�j����	��h	=.�p�}\d�E��4\��pQ��(友�pQ�����pQ���
�S4(}Gz�����Pz��!���Pz�	�A���Pz�
�a���P���>�ņq����5���n}�V��}�[�m|�Dty��_�:����]��+_xɏ������/y�<|��~�����p�������� �?������Cp_���қ�?��WZ��p��d+�_�v?}}���\��뻇�/|���>l����g�����v���}��?����a���}��j���u���=|�������"��X�\�=lw>�'��}L�cT����=嚏1������Ӷ���+Y�i����e�SMM��*�:��8����6Q�IoV;���m���h��o����}R����apC�y{�F�rA�?-q�M��;�ĥÒ�×������C�����?y�n���&�w_�Ň4�$��_~�kv|R�t�V��||����ݔ�ܖ%�eQ��L�)��
����K��(�*����i�Φ.�]ۏS*�zLJ9�ypSdِ,�?��$S'��6-l�V�����SN��wQ������'y���MYܺ��_q�6m�̙4��$�3��6�I�`�Rd�sv�Q7J�����ƦC���{�Gq�$;]�N���%t�$�N�d����j��{�Ĝ,q�ɒ"��^����=�9�_f�lG�����vyyf���vٙ��3����!�YV��e���3ۥg��g�3��w��2�z�RU��ѯ1*�,��C�j�iUj�M[��0Yٹ��?
J����ʦ�شJ���u�3�*Q��An8�)pҏK�xP�qI���Ө������$��/�n�<f��r�M�3�c��iBU���M�'M֕IѓM��۟�n�<+Ma�"���G$�&�� .K�A��#7=~�>�2T��ra<]����y�jrK��㾗g�Ǐ�Yt��lz��	�Iu<�8~��IՔ�����#�U��O�}��d���I��~��w�}��\R��"։�Ǐ>ʟ|�����f��/�Y�w���=��o��l�����F���7���~���lw�;=�a��<��?�ÿ�?�y��כ��|�K����5tV�/�ͳ?/=�>��������t��>3��j�J'h��>�c}��_����';{[�*���HM^�7�m겊�3Uj���s�r~��{���%-5.q]������.-rk�3_�5�կv0��������O���o��������W�?����������-�OWݦ�2%U�����؏��"O�������C4�Q���!���}��篿��??��?�?�_�Ls�5���ad�<-��m~[:ʝu��YQHȨ'FG��~�����������}��_��������Uϔ|���L3���I7�,oG����dee��ٿ���_7�c���qH�沲�D|%�L�H�t�]�t��3$��H3�I�ɨ��c�^�$���Χ��W�ۧ6<��?�(���O�����Ϻ�UQ����xժ�n�"�_�k��_���z�k����o�����o��������P���W�PoV�ެ��嗼���_'�?��_�â�gyb�};!%��1H�럾C�z�/�h�ﶾ|Շw���o޼Y��,_�����������������ǫ�k����8����ji6��pc��joy���g�ˬ�������VV�w?��"S̊'��Y��A���x�Z�fQY�6�UgL�!��:�K�9���:�W�-���}��{}�Z�E��p�齾�7�Z�g���Z0A�4+����A��������T�y��,�XM�|7�c����������mn�<�5���N'Oa�X-�쵨��M�昻��-@������YAn��F�ɓ]��J���nM���� �<�����ik6y"�n��b+O�w���qs5n��Y7����t���y�[��O�����Ůf�tr��i�L{�
�ҩ���.�\��8=^��d�/�W+�W���籫��d\�L�".Ֆ���z@Ob��#�xT�Il�vi"�Ȇ��fb-k��JGW��V��Du���Ny��'�:�KS�^� 7kY�)M�5�Ŏ~�Nd�lٱW&�Xd��]�>i���L�<�d'W�F'���f.Kg���#�`�<�-�E�����z~V�L~�V�̉�'��ufn���OOMk��<�Gd��<�����tk���(��3s�j����UZ@��8s�	���~	���H��h5r�����"��9�t[ ���l~\i��1Z����ɼ��Ş_�5��90?�w��`�q�}�<�~�V�icd�kV��E�d��8瞖�qC���t���(��h5���B�P�j�e�z�a�ͨ4�5�������I�ُ7+M�fZ��o蘱O[\���V���>�gԟ���&M�e��^p��9�ץ�7��}0��_炇�8�{j�<4^����h<؍Z�7;a/��{�+
�
��Ҋ�G\�������� ��J�g"c�|��� fi�V����*��U��iET��jTMg�x��LU�3ۻ�����C���w�b�0����گ���ݟw?�>t?>�^\���PK   �WW��?�(  �            ��    cirkitFile.jsonPK      =   �(    